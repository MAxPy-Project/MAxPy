module adder4(A, B, SUM); 
input  [3:0] A; 
input  [3:0] B; 
output [3:0] SUM;
assign SUM = A + B; 
endmodule
